library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library work;
use work.all;


entity INIT_RAM is
	port(
			clk : in std_logic;
			rst : in std_logic;
			address : in std_logic_vector(8 downto 0);
			data : out std_logic_vector(15 downto 0);
			finished : out std_logic
	);
end INIT_RAM;

architecture INIT_RAM_ARCH of INIT_RAM is

begin

	process(clk, rst)
	begin
	
		if( rst = '1' ) then
			data <= x"0000";
			finished <= '0';
		elsif(clk = '1' and clk'event) then
			finished <= '0';
			case(address) is
			--JPEG Init
			  when '0' & x"00" =>
					data <= x"ff00";
			  when '0' & x"01" =>
					data <= x"2cff";
			  when '0' & x"02" =>
					data <= x"2edf"; -- df
			  when '0' & x"03" =>
					data <= x"ff01";
			  when '0' & x"04" =>
					data <= x"3c32";
			  when '0' & x"05" =>
					data <= x"1100";	
			  when '0' & x"06" =>
					data <= x"0902";
			  when '0' & x"07" =>
					data <= x"0428"; --28
			  when '0' & x"08" =>
					data <= x"13e5";
			  when '0' & x"09" =>
					data <= x"1448";
			  when '0' & x"0A" =>
					data <= x"2c0c";
			  when '0' & x"0B" =>
					data <= x"3378";
			  when '0' & x"0C" =>
					data <= x"3a33";
			  when '0' & x"0D" =>
					data <= x"3bfB";
			  when '0' & x"0E" =>
					data <= x"3e00";
			  when '0' & x"0F" =>
					data <= x"4311";
			  when '0' & x"10" =>
					data <= x"1610";
			  when '0' & x"11" =>
					data <= x"3992";
			  when '0' & x"12" =>
					data <= x"35da";
			  when '0' & x"13" =>
					data <= x"221a";
			  when '0' & x"14" =>
					data <= x"37c3";
			  when '0' & x"15" =>
					data <= x"2300";
			  when '0' & x"16" =>
					data <= x"34c0";
			  when '0' & x"17" =>
					data <= x"361a";
			  when '0' & x"18" =>
					data <= x"0688";
			  when '0' & x"19" =>
					data <= x"07c0";
			  when '0' & x"1A" =>
					data <= x"0d87";
			  when '0' & x"1B" =>
					data <= x"0e41";
			  when '0' & x"1C" =>
					data <= x"4c00";
			  when '0' & x"1D" =>
					data <= x"4800";
			  when '0' & x"1E" =>
					data <= x"5B00";
			  when '0' & x"1F" =>
					data <= x"4203";
			  when '0' & x"20" =>
					data <= x"4a81";
			  when '0' & x"21" =>
					data <= x"2199";
			  when '0' & x"22" =>
					data <= x"2440";
			  when '0' & x"23" =>
					data <= x"2538";
			  when '0' & x"24" =>
					data <= x"2682";
			  when '0' & x"25" =>
					data <= x"5c00";
			  when '0' & x"26" =>
					data <= x"6300";
			  when '0' & x"27" =>
					data <= x"6170";
			  when '0' & x"28" =>
					data <= x"6280";
			  when '0' & x"29" =>
					data <= x"7c05";
			  when '0' & x"2A" =>
					data <= x"2080";
			  when '0' & x"2B" =>
					data <= x"2830";
			  when '0' & x"2C" =>
					data <= x"6c00";
			  when '0' & x"2D" =>
					data <= x"6d80";
			  when '0' & x"2E" =>
					data <= x"6e00";
			  when '0' & x"2F" =>
					data <= x"7002";
			  when '0' & x"30" =>
					data <= x"7194";
			  when '0' & x"31" =>
					data <= x"73c1";
			  when '0' & x"32" =>
					data <= x"1240";
			  when '0' & x"33" =>
					data <= x"1711"; -- 11
			  when '0' & x"34" =>
					data <= x"1843";
			  when '0' & x"35" =>
					data <= x"1900";
			  when '0' & x"36" =>
					data <= x"1a4b";
			  when '0' & x"37" =>
					data <= x"3209"; -- 09
			  when '0' & x"38" =>
					data <= x"37c0";
			  when '0' & x"39" =>
					data <= x"4f60";
			  when '0' & x"3A" =>
					data <= x"50a8";
			  when '0' & x"3B" =>
					data <= x"6d00";
			  when '0' & x"3C" =>
					data <= x"3d38";
			  when '0' & x"3D" =>
					data <= x"463f";
			  when '0' & x"3E" =>
					data <= x"4f60";
			  when '0' & x"3F" =>
					data <= x"0c3c";
			  when '0' & x"40" =>
					data <= x"ff00";
			  when '0' & x"41" =>
					data <= x"e57f";
			  when '0' & x"42" =>
					data <= x"f9c0";
			  when '0' & x"43" =>
					data <= x"4124";
			  when '0' & x"44" =>
					data <= x"e014";
			  when '0' & x"45" =>
					data <= x"76ff";
			  when '0' & x"46" =>
					data <= x"33a0";
			  when '0' & x"47" =>
					data <= x"4220";
			  when '0' & x"48" =>
					data <= x"4318";
			  when '0' & x"49" =>
					data <= x"4c00";
			  when '0' & x"4A" =>
					data <= x"87d5";
			  when '0' & x"4B" =>
					data <= x"883f";
			  when '0' & x"4C" =>
					data <= x"d703";
			  when '0' & x"4D" =>
					data <= x"d910";
			  when '0' & x"4E" =>
					data <= x"d382";
			  when '0' & x"4F" =>
					data <= x"c808";
			  when '0' & x"50" =>
					data <= x"c980";
			  when '0' & x"51" =>
					data <= x"7c00";
			  when '0' & x"52" =>
					data <= x"7d00";
			  when '0' & x"53" =>
					data <= x"7c03";
			  when '0' & x"54" =>
					data <= x"7d48";
			  when '0' & x"55" =>
					data <= x"7d48";
			  when '0' & x"56" =>
					data <= x"7c08";
			  when '0' & x"57" =>
					data <= x"7d20";
			  when '0' & x"58" =>
					data <= x"7d10";
			  when '0' & x"59" =>
					data <= x"7d0e";
			  when '0' & x"5A" =>
					data <= x"9000";
			  when '0' & x"5B" =>
					data <= x"910e";
			  when '0' & x"5C" =>
					data <= x"911a";
			  when '0' & x"5D" =>
					data <= x"9131";
			  when '0' & x"5E" =>
					data <= x"915a";
			  when '0' & x"5F" =>
					data <= x"9169";
			  when '0' & x"60" =>
					data <= x"9175";
			  when '0' & x"61" =>
					data <= x"917e";
			  when '0' & x"62" =>
					data <= x"9188";
			  when '0' & x"63" =>
					data <= x"918f";
			  when '0' & x"64" =>
					data <= x"9196";
			  when '0' & x"65" =>
					data <= x"91a3";
			  when '0' & x"66" =>
					data <= x"91af";
			  when '0' & x"67" =>
					data <= x"91c4";
			  when '0' & x"68" =>
					data <= x"91d7";
			  when '0' & x"69" =>
					data <= x"91e8";
			  when '0' & x"6A" =>
					data <= x"9120";
			  when '0' & x"6B" =>
					data <= x"9200";
			  when '0' & x"6C" =>
					data <= x"9306";
			  when '0' & x"6D" =>
					data <= x"93e3";
			  when '0' & x"6E" =>
					data <= x"9305";
			  when '0' & x"6F" =>
					data <= x"9305";
			  when '0' & x"70" =>
					data <= x"9300";
			  when '0' & x"71" =>
					data <= x"9304";
			  when '0' & x"72" =>
					data <= x"9300";
			  when '0' & x"73" =>
					data <= x"9300";
			  when '0' & x"74" =>
					data <= x"9300";
			  when '0' & x"75" =>
					data <= x"9300";
			  when '0' & x"76" =>
					data <= x"9300";
			  when '0' & x"77" =>
					data <= x"9300";
			  when '0' & x"78" =>
					data <= x"9300";
			  when '0' & x"79" =>
					data <= x"9600";
			  when '0' & x"7A" =>
					data <= x"9708";
			  when '0' & x"7B" =>
					data <= x"9719";
			  when '0' & x"7C" =>
					data <= x"9702";
			  when '0' & x"7D" =>
					data <= x"970c";
			  when '0' & x"7E" =>
					data <= x"9724";
			  when '0' & x"7F" =>
					data <= x"9730";
			  when '0' & x"80" =>
					data <= x"9728";
			  when '0' & x"81" =>
					data <= x"9726";
			  when '0' & x"82" =>
					data <= x"9702";
			  when '0' & x"83" =>
					data <= x"9798";
			  when '0' & x"84" =>
					data <= x"9780";
			  when '0' & x"85" =>
					data <= x"9700";
			  when '0' & x"86" =>
					data <= x"9700";
			  when '0' & x"87" =>
					data <= x"c3ed";
			  when '0' & x"88" =>
					data <= x"a400";
			  when '0' & x"89" =>
					data <= x"a800";
			  when '0' & x"8A" =>
					data <= x"c511";
			  when '0' & x"8B" =>
					data <= x"c651";
			  when '0' & x"8C" =>
					data <= x"bf80";
			  when '0' & x"8D" =>
					data <= x"c710";
			  when '0' & x"8E" =>
					data <= x"b666";
			  when '0' & x"8F" =>
					data <= x"b8A5";
			  when '0' & x"90" =>
					data <= x"b764";
			  when '0' & x"91" =>
					data <= x"b97C";
			  when '0' & x"92" =>
					data <= x"b3af";
			  when '0' & x"93" =>
					data <= x"b497";
			  when '0' & x"94" =>
					data <= x"b5FF";
			  when '0' & x"95" =>
					data <= x"b0C5";
			  when '0' & x"96" =>
					data <= x"b194";
			  when '0' & x"97" =>
					data <= x"b20f";
			  when '0' & x"98" =>
					data <= x"c45c";
			  when '0' & x"99" =>
					data <= x"c064";
			  when '0' & x"9A" =>
					data <= x"c14B";
			  when '0' & x"9B" =>
					data <= x"8c00";
			  when '0' & x"9C" =>
					data <= x"863D";
			  when '0' & x"9D" =>
					data <= x"5000";
			  when '0' & x"9E" =>
					data <= x"51C8";
			  when '0' & x"9F" =>
					data <= x"5296";
			  when '0' & x"A0" =>
					data <= x"5300";
			  when '0' & x"A1" =>
					data <= x"5400";
			  when '0' & x"A2" =>
					data <= x"5500";
			  when '0' & x"A3" =>
					data <= x"5aC8";
			  when '0' & x"A4" =>
					data <= x"5b96";
			  when '0' & x"A5" =>
					data <= x"5c00";
			  when '0' & x"A6" =>
					data <= x"d300";	--//when '0' & x"A0" =>data <= x"d37f";
			  when '0' & x"A7" =>
					data <= x"c3ed";
			  when '0' & x"A8" =>
					data <= x"7f00";
			  when '0' & x"A9" =>
					data <= x"da00";
			  when '0' & x"AA" =>
					data <= x"e51f";
			  when '0' & x"AB" =>
					data <= x"e167";
			  when '0' & x"AC" =>
					data <= x"e000";
			  when '0' & x"AD" =>
					data <= x"dd7f";
			  when '0' & x"AE" =>
					data <= x"0500";
			  when '0' & x"AF" =>
					data <= x"1240";
			  when '0' & x"B0" =>
					data <= x"d304";	--//when '0' & x"B0" =>data <= x"d37f";
			  when '0' & x"B1" =>
					data <= x"c016";
			  when '0' & x"B2" =>
					data <= x"C112";
			  when '0' & x"B3" =>
					data <= x"8c00";
			  when '0' & x"B4" =>
					data <= x"863d";
			  when '0' & x"B5" =>
					data <= x"5000";
			  when '0' & x"B6" =>
					data <= x"512C";
			  when '0' & x"B7" =>
					data <= x"5224";
			  when '0' & x"B8" =>
					data <= x"5300";
			  when '0' & x"B9" =>
					data <= x"5400";
			  when '0' & x"BA" =>
					data <= x"5500";
			  when '0' & x"BB" =>
					data <= x"5A2c";
			  when '0' & x"BC" =>
					data <= x"5b24";
			  when '0' & x"BD" =>
					data <= x"5c00";
			  when '0' & x"BE" =>
					data <= x"FF00";
			  when '0' & x"BF" =>
					data <= x"0500";
			  when '0' & x"C0" =>
					data <= x"DA10";
			  when '0' & x"C1" =>
					data <= x"D703";
			  when '0' & x"C2" =>
					data <= x"DF00";
			  when '0' & x"C3" =>
					data <= x"3380";
			  when '0' & x"C4" =>
					data <= x"3C40";
			  when '0' & x"C5" =>
					data <= x"e177";
			  when '0' & x"C6" =>
					data <= x"0000";
			  -- From YUV422 Mode
			  when '0' & x"C7" =>
					data <= x"FF00";
			  when '0' & x"C8" =>
					data <= x"0500";
			  when '0' & x"C9" =>
					data <= x"DA10";
			  when '0' & x"CA" =>
					data <= x"D703";
			  when '0' & x"CB" =>
					data <= x"DF00";
			  when '0' & x"CC" =>
					data <= x"3380";
			  when '0' & x"CD" =>
					data <= x"3C40";
			  when '0' & x"CE" =>
					data <= x"e177";
			  when '0' & x"CF" =>
					data <= x"0000"; 
				-- More Jpeg Stuff
			  when '0' & x"D0" =>
					data <= x"e014";
			  when '0' & x"D1" =>
					data <= x"e177";
			  when '0' & x"D2" =>
					data <= x"e51f";
			  when '0' & x"D3" =>
					data <= x"d703";
			  when '0' & x"D4" =>
					data <= x"da10"; -- 10
			  when '0' & x"D5" =>
					data <= x"e000";
			  when '0' & x"D6" =>
					data <= x"FF01";
			  when '0' & x"D7" =>
					data <= x"0408";
			 --800 x 600 jpeG
				when '0' & x"D8" =>
					data <= x"ff01";
			   when '0' & x"D9" =>
					data <= x"1100";
				when '0' & x"DA" =>
					data <= x"1240"; --// Bit[6:4]: Resolution selection//0x02为彩条
				when '0' & x"DB" =>
					data <= x"1711"; -- 11
				when '0' & x"DC" =>
					data <= x"1843"; --75 to 43
				when '0' & x"DD" =>
					data <= x"3209"; --36 to 09
				when '0' & x"DE" =>
					data <= x"1900"; -- 01 to 00
				when '0' & x"DF" =>
					data <= x"1a4b"; -- 94 to 4b
				when '0' & x"E0" =>
					data <= x"030A"; -- 0F to 0A
				when '0' & x"E1" =>
					data <= x"3740"; -- unknown
				when '0' & x"E2" =>
					data <= x"4fbb"; 
				when '0' & x"E3" =>
					data <= x"509c";
				when '0' & x"E4" =>
					data <= x"5a57";
				when '0' & x"E5" =>
					data <= x"6d80";
				when '0' & x"E6" =>
					data <= x"3d34";
				when '0' & x"E7" =>
					data <= x"3902";
				when '0' & x"E8" =>
					data <= x"3588";
				when '0' & x"E9" =>
					data <= x"220a";
				when '0' & x"EA" =>
					data <= x"3740";
				when '0' & x"EB" =>
					data <= x"34a0";
				when '0' & x"EC" =>
					data <= x"0602";
				when '0' & x"ED" =>
					data <= x"0db7";
				when '0' & x"EE" =>
					data <= x"0e01";		
				when '0' & x"EF" =>
					data <= x"ff00";
				when '0' & x"F0" =>
					data <= x"e004";
				when '0' & x"F1" =>
					data <= x"c064"; -- c8 to 64
				when '0' & x"F2" =>
					data <= x"c14b"; -- 96 to 4b
				when '0' & x"F3" =>
					data <= x"8635";
				when '0' & x"F4" =>
					data <= x"5080"; -- 89 to 80
				when '0' & x"F5" =>
					data <= x"51c8"; -- 90 to c8
				when '0' & x"F6" => 
					data <= x"5296"; -- 2c to 96
				when '0' & x"F7" =>
					data <= x"5300"; -- 00
				when '0' & x"F8" =>
					data <= x"5400"; -- 00
				when '0' & x"F9" =>
					data <= x"5500"; -- 88 to 00
				when '0' & x"FA" =>
					data <= x"5700"; -- 00
				when '0' & x"FB" =>
					data <= x"5ac8"; -- c8
				when '0' & x"FC" =>
					data <= x"5b96"; -- 96
				when '0' & x"FD" =>
					data <= x"5c00"; -- 00
				when '0' & x"FE" =>
					data <= x"d302"; 
				when '0' & x"FF" =>
					data <= x"e000"; -- 00				 
				when '1' & x"00" =>
					data <= x"ff01";
				-- Custom 
				when '1' & x"01" =>
					data <= x"1140"; -- 00 MASTER -- 40 SLAVE
				when '1' & x"02" =>
					data <= x"0906"; -- 06 SLV MODE -- 02 MASTER
				when '1' & x"03" =>
					data <= x"1248"; -- 48 -- SVGA MASTER MODE
				-- MASTER SVGA ESTABLISHED.
				-- TIMINGS :-

			
			
			
			

			
			
				when others =>
					data <= x"0000";
					finished <= '1';
					
				
			
					
					
				end case;
		end if;
	end process;

end INIT_RAM_ARCH;