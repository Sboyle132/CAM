library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library work;
use work.all;


entity INIT_RAM is
	port(
			clk : in std_logic;
			rst : in std_logic;
			address : in std_logic_vector(8 downto 0);
			data : out std_logic_vector(15 downto 0);
			finished : out std_logic
	);
end INIT_RAM;

architecture INIT_RAM_ARCH of INIT_RAM is

begin

	process(clk, rst)
	begin
	
		if( rst = '1' ) then
			data <= x"0000";
			finished <= '0';
		elsif(clk = '1' and clk'event) then
			finished <= '0';
			case(address) is
			when '0' & x"00" =>
				data <= x"ff01";
			when '0' & x"01" =>
				data <= x"1280";
			when '0' & x"02" =>
				data <= x"ff00";
			when '0' & x"03" =>
				data <= x"2cff";
			when '0' & x"04" =>
				data <= x"2edf";
			when '0' & x"05" =>
				data <= x"ff01";
			when '0' & x"06" =>
				data <= x"3c32";
			when '0' & x"07" =>
				data <= x"1101"; -- 01 MASTER -- 41 SLAVE
			when '0' & x"08" =>
				data <= x"0902"; -- 06 SLV MODE -- 02 MASTER
			when '0' & x"09" =>
				data <= x"0428";
			when '0' & x"0A" =>
				data <= x"13e5";
			when '0' & x"0B" =>
				data <= x"1448";
			when '0' & x"0C" =>
				data <= x"2c0c";
			when '0' & x"0D" =>
				data <= x"3378";
			when '0' & x"0E" =>
				data <= x"3a33";
			when '0' & x"0F" =>
				data <= x"3bfB";
			when '0' & x"10" =>
				data <= x"3e00";
			when '0' & x"11" =>
				data <= x"4311";
			when '0' & x"12" =>
				data <= x"1610";
			when '0' & x"13" =>
				data <= x"3992";
			when '0' & x"14" =>
				data <= x"35da";
			when '0' & x"15" =>
				data <= x"221a";
			when '0' & x"16" =>
				data <= x"37c3";
			when '0' & x"17" =>
				data <= x"2300";
			when '0' & x"18" =>
				data <= x"34c0";
			when '0' & x"19" =>
				data <= x"361a";
			when '0' & x"1A" =>
				data <= x"0688";
			when '0' & x"1B" =>
				data <= x"07c0";
			when '0' & x"1C" =>
				data <= x"0d87";
			when '0' & x"1D" =>
				data <= x"0e41";
			when '0' & x"1E" =>
				data <= x"4c00";
			when '0' & x"1F" =>
				data <= x"4800";
			when '0' & x"20" =>
				data <= x"5B00";
			when '0' & x"21" =>
				data <= x"4203";
			when '0' & x"22" =>
				data <= x"4a81";
			when '0' & x"23" =>
				data <= x"2199";
			when '0' & x"24" =>
				data <= x"2440";
			when '0' & x"25" =>
				data <= x"2538";
			when '0' & x"26" =>
				data <= x"2682";
			when '0' & x"27" =>
				data <= x"5c00";
			when '0' & x"28" =>
				data <= x"6300";
			when '0' & x"29" =>
				data <= x"6170";
			when '0' & x"2A" =>
				data <= x"6280";
			when '0' & x"2B" =>
				data <= x"7c05";
			when '0' & x"2C" =>
				data <= x"2080";
			when '0' & x"2D" =>
				data <= x"2830";
			when '0' & x"2E" =>
				data <= x"6c00";
			when '0' & x"2F" =>
				data <= x"6d80";
			when '0' & x"30" =>
				data <= x"6e00";
			when '0' & x"31" =>
				data <= x"7002";
			when '0' & x"32" =>
				data <= x"7194";
			when '0' & x"33" =>
				data <= x"73c1";
			when '0' & x"34" =>
				data <= x"1240"; -- 40 MASTER MODE -- 48 SLAVE MODE
			when '0' & x"35" =>
				data <= x"1711";
			when '0' & x"36" =>
				data <= x"1843";
			when '0' & x"37" =>
				data <= x"1900";
			when '0' & x"38" =>
				data <= x"1a4b";
			when '0' & x"39" =>
				data <= x"3209";
			when '0' & x"3A" =>
				data <= x"37c0";
			when '0' & x"3B" =>
				data <= x"4f60";
			when '0' & x"3C" =>
				data <= x"50a8";
			when '0' & x"3D" =>
				data <= x"6d00";
			when '0' & x"3E" =>
				data <= x"3d38";
			when '0' & x"3F" =>
				data <= x"463f";
			when '0' & x"40" =>
				data <= x"4f60";
			when '0' & x"41" =>
				data <= x"0c3c";
			when '0' & x"42" =>
				data <= x"ff00";
			when '0' & x"43" =>
				data <= x"e57f";
			when '0' & x"44" =>
				data <= x"f9c0";
			when '0' & x"45" =>
				data <= x"4124";
			when '0' & x"46" =>
				data <= x"e014";
			when '0' & x"47" =>
				data <= x"76ff";
			when '0' & x"48" =>
				data <= x"33a0";
			when '0' & x"49" =>
				data <= x"4220";
			when '0' & x"4A" =>
				data <= x"4318";
			when '0' & x"4B" =>
				data <= x"4c00";
			when '0' & x"4C" =>
				data <= x"87d5";
			when '0' & x"4D" =>
				data <= x"883f";
			when '0' & x"4E" =>
				data <= x"d703";
			when '0' & x"4F" =>
				data <= x"d910";
			when '0' & x"50" =>
				data <= x"d382";
			when '0' & x"51" =>
				data <= x"c808";
			when '0' & x"52" =>
				data <= x"c980";
			when '0' & x"53" =>
				data <= x"7c00";
			when '0' & x"54" =>
				data <= x"7d00";
			when '0' & x"55" =>
				data <= x"7c03";
			when '0' & x"56" =>
				data <= x"7d48";
			when '0' & x"57" =>
				data <= x"7d48";
			when '0' & x"58" =>
				data <= x"7c08";
			when '0' & x"59" =>
				data <= x"7d20";
			when '0' & x"5A" =>
				data <= x"7d10";
			when '0' & x"5B" =>
				data <= x"7d0e";
			when '0' & x"5C" =>
				data <= x"9000";
			when '0' & x"5D" =>
				data <= x"910e";
			when '0' & x"5E" =>
				data <= x"911a";
			when '0' & x"5F" =>
				data <= x"9131";
			when '0' & x"60" =>
				data <= x"915a";
			when '0' & x"61" =>
				data <= x"9169";
			when '0' & x"62" =>
				data <= x"9175";
			when '0' & x"63" =>
				data <= x"917e";
			when '0' & x"64" =>
				data <= x"9188";
			when '0' & x"65" =>
				data <= x"918f";
			when '0' & x"66" =>
				data <= x"9196";
			when '0' & x"67" =>
				data <= x"91a3";
			when '0' & x"68" =>
				data <= x"91af";
			when '0' & x"69" =>
				data <= x"91c4";
			when '0' & x"6A" =>
				data <= x"91d7";
			when '0' & x"6B" =>
				data <= x"91e8";
			when '0' & x"6C" =>
				data <= x"9120";
			when '0' & x"6D" =>
				data <= x"9200";
			when '0' & x"6E" =>
				data <= x"9306";
			when '0' & x"6F" =>
				data <= x"93e3";
			when '0' & x"70" =>
				data <= x"9305";
			when '0' & x"71" =>
				data <= x"9305";
			when '0' & x"72" =>
				data <= x"9300";
			when '0' & x"73" =>
				data <= x"9304";
			when '0' & x"74" =>
				data <= x"9300";
			when '0' & x"75" =>
				data <= x"9300";
			when '0' & x"76" =>
				data <= x"9300";
			when '0' & x"77" =>
				data <= x"9300";
			when '0' & x"78" =>
				data <= x"9300";
			when '0' & x"79" =>
				data <= x"9300";
			when '0' & x"7A" =>
				data <= x"9300";
			when '0' & x"7B" =>
				data <= x"9600";
			when '0' & x"7C" =>
				data <= x"9708";
			when '0' & x"7D" =>
				data <= x"9719";
			when '0' & x"7E" =>
				data <= x"9702";
			when '0' & x"7F" =>
				data <= x"970c";
			when '0' & x"80" =>
				data <= x"9724";
			when '0' & x"81" =>
				data <= x"9730";
			when '0' & x"82" =>
				data <= x"9728";
			when '0' & x"83" =>
				data <= x"9726";
			when '0' & x"84" =>
				data <= x"9702";
			when '0' & x"85" =>
				data <= x"9798";
			when '0' & x"86" =>
				data <= x"9780";
			when '0' & x"87" =>
				data <= x"9700";
			when '0' & x"88" =>
				data <= x"9700";
			when '0' & x"89" =>
				data <= x"c3ed";
			when '0' & x"8A" =>
				data <= x"a400";
			when '0' & x"8B" =>
				data <= x"a800";
			when '0' & x"8C" =>
				data <= x"c511";
			when '0' & x"8D" =>
				data <= x"c651";
			when '0' & x"8E" =>
				data <= x"bf80";
			when '0' & x"8F" =>
				data <= x"c710";
			when '0' & x"90" =>
				data <= x"b666";
			when '0' & x"91" =>
				data <= x"b8A5";
			when '0' & x"92" =>
				data <= x"b764";
			when '0' & x"93" =>
				data <= x"b97C";
			when '0' & x"94" =>
				data <= x"b3af";
			when '0' & x"95" =>
				data <= x"b497";
			when '0' & x"96" =>
				data <= x"b5FF";
			when '0' & x"97" =>
				data <= x"b0C5";
			when '0' & x"98" =>
				data <= x"b194";
			when '0' & x"99" =>
				data <= x"b20f";
			when '0' & x"9A" =>
				data <= x"c45c";
			when '0' & x"9B" =>
				data <= x"c064";
			when '0' & x"9C" =>
				data <= x"c14B";
			when '0' & x"9D" =>
				data <= x"8c00";
			when '0' & x"9E" =>
				data <= x"863D";
			when '0' & x"9F" =>
				data <= x"5000";
			when '0' & x"A0" =>
				data <= x"51C8";
			when '0' & x"A1" =>
				data <= x"5296";
			when '0' & x"A2" =>
				data <= x"5300";
			when '0' & x"A3" =>
				data <= x"5400";
			when '0' & x"A4" =>
				data <= x"5500";
			when '0' & x"A5" =>
				data <= x"5aC8";
			when '0' & x"A6" =>
				data <= x"5b96";
			when '0' & x"A7" =>
				data <= x"5c00";
			when '0' & x"A8" =>
				data <= x"d382";
			when '0' & x"A9" =>
				data <= x"c3ed";
			when '0' & x"AA" =>
				data <= x"7f00";
			when '0' & x"AB" =>
				data <= x"da00";
			when '0' & x"AC" =>
				data <= x"e51f";
			when '0' & x"AD" =>
				data <= x"e167";
			when '0' & x"AE" =>
				data <= x"e000";
			when '0' & x"AF" =>
				data <= x"dd7f";
			when '0' & x"B0" =>
				data <= x"0500";
			when '0' & x"B1" =>
				data <= x"ff01";
	
	













	
	
	
--				when '0' & x"00" =>
--					data <= x"ff01";
--				when '0' & x"01" =>
--					data <= x"ff01";
--				when '0' & x"02" =>
--					data <= x"2cff";
--				when '0' & x"03" =>
--					data <= x"2edf";
--				when '0' & x"04" =>
--					data <= x"ff01";
--				when '0' & x"05" =>	
--					data <= x"3c32";
--				when '0' & x"06" =>
--					data <= x"1101";
--				when '0' & x"07" =>
--					data <= x"0902";
--				when '0' & x"08" =>
--					data <= x"0428";
--				when '0' & x"09" =>
--					data <= x"13e5";
--				when '0' & x"0A" =>
--					data <= x"1448";
--				when '0' & x"0B" =>
--					data <= x"2c0c";
--				when '0' & x"0C" =>
--					data <= x"3378";
--				when '0' & x"0D" =>
--					data <= x"3a33";  
-- 				when '0' & x"0E" =>
--					data <= x"3bfb";  
-- 				when '0' & x"0F" =>
--					data <= x"3e00";  
-- 				when '0' & x"10" =>
--					data <= x"4311";  
-- 				when '0' & x"11" =>
--					data <= x"1610";  
-- 				when '0' & x"12" =>
--					data <= x"3992";  
-- 				when '0' & x"13" =>
--					data <= x"35DA";  
-- 				when '0' & x"14" =>
--					data <= x"221A";  
-- 				when '0' & x"15" =>
--					data <= x"37C3";  
-- 				when '0' & x"16" =>
--					data <= x"2300";  
-- 				when '0' & x"17" =>
--					data <= x"34C0";  
-- 				when '0' & x"18" =>
--					data <= x"0602";
--		
-- 				when '0' & x"19" =>
--					data <= x"0688";  
-- 				when '0' & x"1A" =>
--					data <= x"07c0";  
-- 				when '0' & x"1B" =>
--					data <= x"0D87";  
-- 				when '0' & x"1C" =>
--					data <= x"0E41";  
-- 				when '0' & x"1D" =>
--					data <= x"4C00";  
-- 				when '0' & x"1E" =>
--					data <= x"4a81";
-- 				when '0' & x"1F" =>
--					 data <= x"2199";  
-- 				when '0' & x"20" =>
--					data <= x"2199";  		
-- 				when '0' & x"21" =>
--					data <= x"2538";
-- 				when '0' & x"22" =>
--					data <= x"2682";
-- 				when '0' & x"23" =>
--					data <= x"5c00";
-- 				when '0' & x"24" =>
--					data <= x"6300";
-- 				when '0' & x"25" =>
--					data <= x"4622";
-- 				when '0' & x"26" =>
--					data <= x"0c3a";  
-- 				when '0' & x"27" =>
--					data <= x"5d55";
-- 				when '0' & x"28" =>
--					data <= x"5e7d";  
-- 				when '0' & x"29" =>
--					data <= x"5f7d";  
-- 				when '0' & x"2A" =>
--					data <= x"6055";  
-- 				when '0' & x"2B" =>
--					data <= x"6170";  
-- 				when '0' & x"2C" =>
--					data <= x"6280";  
-- 				when '0' & x"2D" =>
--					data <= x"7c05";  
-- 				when '0' & x"2E" =>
--					data <= x"2080";  
-- 				when '0' & x"2F" => 
--					data <= x"2830";  
-- 				when '0' & x"30" =>
--					data <= x"6c00";  
-- 				when '0' & x"31" =>
--					data <= x"6d80";  
-- 				when '0' & x"32" =>
--					data <= x"6e00";  
-- 				when '0' & x"33" =>
--					data <= x"7002";  
-- 				when '0' & x"34" =>
--					data <= x"7194";  
-- 				when '0' & x"35" =>
--					data <= x"73c1";  
-- 				when '0' & x"36" =>
--					data <= x"3d34";  
-- 				when '0' & x"37" =>
--					data <= x"1204";  
-- 				when '0' & x"38" =>
--					data <= x"5a57";  
-- 				when '0' & x"39" =>
--					data <= x"4fbb";  
-- 				when '0' & x"3A" =>
--					data <= x"509c";  
-- 				when '0' & x"3B" =>
--					data <= x"ff00";  
-- 				when '0' & x"3C" =>
--					data <= x"e57f";  
-- 				when '0' & x"3D" =>
--					data <= x"f9c0";  
-- 				when '0' & x"3E" =>
--					data <= x"4124";  
-- 				when '0' & x"3F" =>
--					data <= x"e014";  
-- 				when '0' & x"40" =>
--					data <= x"76ff";  
-- 				when '0' & x"41" =>
--					data <= x"33a0";  
-- 				when '0' & x"42" =>
--					data <= x"4220";  
-- 				when '0' & x"43" =>
--					data <= x"4318";  
-- 				when '0' & x"44" =>
--					data <= x"4c00";  
-- 				when '0' & x"45" =>
--					data <= x"87d0";  
-- 				when '0' & x"46" =>
--					data <= x"883f";  
-- 				when '0' & x"47" =>
--					data <= x"d703";  
-- 				when '0' & x"48" =>
--					data <= x"d910";  
-- 				when '0' & x"49" =>
--					data <= x"d382";  
-- 				when '0' & x"4A" =>
--					data <= x"c808";  
-- 				when '0' & x"4B" =>
--					data <= x"c980";  
-- 				when '0' & x"4C" =>
--					data <= x"7c00";  
-- 				when '0' & x"4D" =>
--					data <= x"7d00";  
-- 				when '0' & x"4E" =>
--					data <= x"7c03";  
-- 				when '0' & x"4F" =>
--					data <= x"7d48";  
-- 				when '0' & x"50" =>
--					data <= x"7d48";  
-- 				when '0' & x"51" =>
--					data <= x"7c08";  
-- 				when '0' & x"52" =>
--					data <= x"7d20";  
-- 				when '0' & x"53" =>
--					data <= x"7d10";  
-- 				when '0' & x"54" =>
--					data <= x"7d0e";  
-- 				when '0' & x"55" =>
--					data <= x"9000";  
-- 				when '0' & x"56" =>
--					data <= x"910e";  
-- 				when '0' & x"57" =>
--					data <= x"911a";  
-- 				when '0' & x"58" => 
--					data <= x"9131";  
-- 				when '0' & x"59" =>
--					data <= x"915a";  
-- 				when '0' & x"5A" =>
--					data <= x"9169";  
-- 				when '0' & x"5B" =>
--					data <= x"9175";  
-- 				when '0' & x"5C" =>
--					data <= x"917e";  
-- 				when '0' & x"5D" =>
--					data <= x"9188";  
-- 				when '0' & x"5E" =>
--					data <= x"918f";  
-- 				when '0' & x"5F" => 
--					data <= x"9196";  
-- 				when '0' & x"60" =>
--					data <= x"91a3";  
-- 				when '0' & x"61" =>
--					data <= x"91af";  
-- 				when '0' & x"62" =>
--					data <= x"91c4";  
-- 				when '0' & x"63" =>
--					data <= x"91d7";  
-- 				when '0' & x"64" =>
--					data <= x"91e8";  
-- 				when '0' & x"65" =>
--					data <= x"9120";  
-- 				when '0' & x"66" =>
--					data <= x"9200";  
-- 				when '0' & x"67" =>
--					data <= x"9306";  
-- 				when '0' & x"68" =>
--					data <= x"93e3";  
-- 				when '0' & x"69" =>
--					data <= x"9303";  
-- 				when '0' & x"6A" =>
--					data <= x"9303";  
-- 				when '0' & x"6B" =>
--					data <= x"9300";  
-- 				when '0' & x"6C" =>
--					data <= x"9302";  
-- 				when '0' & x"6D" =>
--					data <= x"9300";  
-- 				when '0' & x"6E" =>
--					data <= x"9300";  
-- 				when '0' & x"6F" =>
--					data <= x"9300";  
-- 				when '0' & x"70" =>
--					data <= x"9300";  
-- 				when '0' & x"71" =>
--					data <= x"9300";  
-- 				when '0' & x"72" =>
--					data <= x"9300";  
-- 				when '0' & x"73" =>
--					data <= x"9300";  
-- 				when '0' & x"74" =>
--					data <= x"9600";  
-- 				when '0' & x"75" =>
--					data <= x"9708";  
-- 				when '0' & x"76" =>
--					data <= x"9719";  
-- 				when '0' & x"77" =>
--					data <= x"9702";  
-- 				when '0' & x"78" =>
--					data <= x"970c";  
-- 				when '0' & x"79" =>
--					data <= x"9724";  
-- 				when '0' & x"7A" =>
--					data <= x"9730";  
-- 				when '0' & x"7B" =>
--					data <= x"9728";  
-- 				when '0' & x"7C" =>
--					data <= x"9726";  
-- 				when '0' & x"7D" =>
--					data <= x"9702";  
-- 				when '0' & x"7E" =>
--					data <= x"9798";  
-- 				when '0' & x"7F" => 
--					data <= x"9780";  
-- 				when '0' & x"80" => 
--					data <= x"9700";  
-- 				when '0' & x"81" => 
--					data <= x"9700";  
-- 				when '0' & x"82" => 
--					data <= x"a400";  
-- 				when '0' & x"83" => 
--					data <= x"a800";  
-- 				when '0' & x"84" => 
--					data <= x"c511";  
-- 				when '0' & x"85" => 
--					data <= x"c651";  
-- 				when '0' & x"86" => 
--					data <= x"bf80";  
-- 				when '0' & x"87" => 
--					data <= x"c710";  
-- 				when '0' & x"88" => 
--					data <= x"b666";  
-- 				when '0' & x"89" => 
--					data <= x"b8a5";  
-- 				when '0' & x"8A" => 
--					data <= x"b764";  
-- 				when '0' & x"8B" => 
--					data <= x"b97c";  
-- 				when '0' & x"8C" => 
--					data <= x"b3af";  
-- 				when '0' & x"8D" => 
--					data <= x"b497";  
-- 				when '0' & x"8E" => 
--					data <= x"b5ff";  
-- 				when '0' & x"8F" => 
--					data <= x"b0c5";  
-- 				when '0' & x"90" => 
--					data <= x"b194";  
-- 				when '0' & x"91" => 
--					data <= x"b20f";  
-- 				when '0' & x"92" => 
--					data <= x"c45c";  
-- 				when '0' & x"93" => 
--					data <= x"a600";  
-- 				when '0' & x"94" => 
--					data <= x"a720";  
-- 				when '0' & x"95" => 
--					data <= x"a7d8";  
-- 				when '0' & x"96" => 
--					data <= x"a71b";  
-- 				when '0' & x"97" => 
--					data <= x"a731";  
-- 				when '0' & x"98" => 
--					data <= x"a700";  
-- 				when '0' & x"99" => 
--					data <= x"a718";  
-- 				when '0' & x"9A" => 
--					data <= x"a720";  
-- 				when '0' & x"9B" => 
--					data <= x"a7d8";  
-- 				when '0' & x"9C" => 
--					data <= x"a719";  
-- 				when '0' & x"9D" => 
--					data <= x"a731";  
-- 				when '0' & x"9E" => 
--					data <= x"a700";  
-- 				when '0' & x"9F" => 
--					data <= x"a718";  
-- 				when '0' & x"A0" => 
--					data <= x"a720";  
-- 				when '0' & x"A1" => 
--					data <= x"a7d8";  
-- 				when '0' & x"A2" => 
--					data <= x"a719";  
-- 				when '0' & x"A3" => 
--					data <= x"a731";  
-- 				when '0' & x"A4" => 
--					data <= x"a700";  
-- 				when '0' & x"A5" => 
--					data <= x"a718";  
-- 				when '0' & x"A6" => 
--					data <= x"7f00";  
-- 				when '0' & x"A7" => 
--					data <= x"e51f";  
-- 				when '0' & x"A8" => 
--					data <= x"e177";  
-- 				when '0' & x"A9" => 
--					data <= x"dd7f";  
-- 				when '0' & x"AA" => 
--					data <= x"c20e";  
-- 				when '0' & x"AB" => 
--					data <= x"ff00";  
-- 				when '0' & x"AC" => 
--					data <= x"e004";  
-- 				when '0' & x"AD" => 
--					data <= x"c0c8";  
-- 				when '0' & x"AE" => 
--					data <= x"c196";  
-- 				when '0' & x"AF" => 
--					data <= x"863d";  
-- 				when '0' & x"B0" => 
--					data <= x"5190";  
-- 				when '0' & x"B1" => 
--					data <= x"522c";  
-- 				when '0' & x"B2" => 
--					data <= x"5300";  
-- 				when '0' & x"B3" => 
--					data <= x"5400";  
-- 				when '0' & x"B4" => 
--					data <= x"5588";  
-- 				when '0' & x"B5" => 
--					data <= x"5700";  
-- 				when '0' & x"B6" => 
--					data <= x"5092";  
-- 				when '0' & x"B7" => 
--					data <= x"5a50";  
-- 				when '0' & x"B8" => 
--					data <= x"5b3c";  
-- 				when '0' & x"B9" => 
--					data <= x"5c00";  
-- 				when '0' & x"BA" => 
--					data <= x"d304";  
-- 				when '0' & x"BB" => 
--					data <= x"e000";  
-- 				when '0' & x"BC" => 
--					data <= x"ff00";  
-- 				when '0' & x"BD" => 
--					data <= x"B500";  
-- 				when '0' & x"BE" =>
--					data <= x"da08";  
-- 				when '0' & x"BF" => 
--					data <= x"d703";  
-- 				when '0' & x"C0" => 
--					data <= x"e000";  
-- 				when '0' & x"C1" => 
--					data <= x"0500";  
-- 				when '0' & x"C2" => 			
--					data <= x"ffff";  			

----------- CONFIG 2
--				when '0' & x"00" =>
--					data <= x"FF01";
--				when '0' & x"01" =>
--					data <= x"1280";
--				when '0' & x"02" =>
--					data <= x"FF00";
--				when '0' & x"03" =>
--					data <= x"2CFF";
--				when '0' & x"04" =>
--					data <= x"2EDF";
--				when '0' & x"05" =>
--					data <= x"FF01";
--				when '0' & x"06" =>
--					data <= x"3C32";
--				when '0' & x"07" =>
--					data <= x"1101";
--				when '0' & x"08" =>
--					data <= x"1101";
--				when '0' & x"09" =>
--					data <= x"0902";
--				when '0' & x"0A" =>
--					data <= x"0420";
--				when '0' & x"0B" =>
--					data <= x"13E5";
--				when '0' & x"0C" =>
--					data <= x"1448";
--				when '0' & x"0D" =>
--					data <= x"2C0C";
--				when '0' & x"0E" =>
--					data <= x"3378";
--				when '0' & x"0F" =>
--					data <= x"3A33";
--				when '0' & x"10" =>
--					data <= x"3BFB";
--				when '0' & x"11" =>
--					data <= x"3E00";
--				when '0' & x"12" =>
--					data <= x"4311";
--				when '0' & x"13" =>
--					data <= x"1610";
--				when '0' & x"14" =>
--					data <= x"3992";
--				when '0' & x"15" =>
--					data <= x"35DA";
--				when '0' & x"16" =>
--					data <= x"221A";
--				when '0' & x"17" =>
--					data <= x"37C3";
--				when '0' & x"18" =>
--					data <= x"2300";
--				when '0' & x"19" =>
--					data <= x"34C0";
--				when '0' & x"1A" =>
--					data <= x"361A";
--				when '0' & x"1B" =>
--					data <= x"0688";
--				when '0' & x"1C" =>
--					data <= x"07C0";
--				when '0' & x"1D" =>
--					data <= x"0D87";
--				when '0' & x"1E" =>
--					data <= x"0E41";
--				when '0' & x"1F" =>
--					data <= x"4C00";
--				when '0' & x"20" =>
--					data <= x"4800";
--				when '0' & x"21" =>
--					data <= x"5B00";
--				when '0' & x"22" =>
--					data <= x"4203";
--				when '0' & x"23" =>
--					data <= x"4A81";
--				when '0' & x"24" =>
--					data <= x"2199";
--				when '0' & x"25" =>
--					data <= x"2440";
--				when '0' & x"26" =>
--					data <= x"2538";
--				when '0' & x"27" =>
--					data <= x"2682";
--				when '0' & x"28" =>
--					data <= x"5C00";
--				when '0' & x"29" =>
--					data <= x"6300";
--				when '0' & x"2A" =>
--					data <= x"4600";
--				when '0' & x"2B" =>
--					data <= x"0C3C";
--				when '0' & x"2C" =>
--					data <= x"6170";
--				when '0' & x"2D" =>
--					data <= x"6280";
--				when '0' & x"2E" =>
--					data <= x"7C05";
--				when '0' & x"2F" =>
--					data <= x"2080";
--				when '0' & x"30" =>
--					data <= x"2830";
--				when '0' & x"31" =>
--					data <= x"6C00";
--				when '0' & x"32" =>
--					data <= x"6D80";
--				when '0' & x"33" =>
--					data <= x"6E00";
--				when '0' & x"34" =>
--					data <= x"7002";
--				when '0' & x"35" =>
--					data <= x"7194";
--				when '0' & x"36" =>
--					data <= x"73C1";
--				when '0' & x"37" =>
--					data <= x"1240";
--				when '0' & x"38" =>
--					data <= x"1711";
--				when '0' & x"39" =>
--					data <= x"1839";
--				when '0' & x"3A" =>
--					data <= x"1900";
--				when '0' & x"3B" =>
--					data <= x"1A3C";
--				when '0' & x"3C" =>
--					data <= x"3209";
--				when '0' & x"3D" =>
--					data <= x"37C0";
--				when '0' & x"3E" =>
--					data <= x"4FCA";
--				when '0' & x"3F" =>
--					data <= x"50A8";
--				when '0' & x"40" =>
--					data <= x"5A23";
--				when '0' & x"41" =>
--					data <= x"6D00";
--				when '0' & x"42" =>
--					data <= x"3D38";
--				when '0' & x"43" =>
--					data <= x"FF00";
--				when '0' & x"44" =>
--					data <= x"E57F";
--				when '0' & x"45" =>
--					data <= x"F9C0";
--				when '0' & x"46" =>
--					data <= x"4124";
--				when '0' & x"47" =>
--					data <= x"E014";
--				when '0' & x"48" =>
--					data <= x"76FF";
--				when '0' & x"49" =>
--					data <= x"33A0";
--				when '0' & x"4A" =>
--					data <= x"4420";
--				when '0' & x"4B" =>
--					data <= x"4318";
--				when '0' & x"4C" =>
--					data <= x"4C00";
--				when '0' & x"4D" =>
--					data <= x"87D5";
--				when '0' & x"4E" =>
--					data <= x"883F";
--				when '0' & x"4F" =>
--					data <= x"D703";
--				when '0' & x"50" =>
--					data <= x"D910";
--				when '0' & x"51" =>
--					data <= x"D382";
--				when '0' & x"52" =>
--					data <= x"C808";
--				when '0' & x"53" =>
--					data <= x"C980";
--				when '0' & x"54" =>
--					data <= x"7C00";
--				when '0' & x"55" =>
--					data <= x"7D00";
--				when '0' & x"56" =>
--					data <= x"7C03";
--				when '0' & x"57" =>
--					data <= x"7D48";
--				when '0' & x"58" =>
--					data <= x"7C08";
--				when '0' & x"59" =>
--					data <= x"7D20";
--				when '0' & x"5A" =>
--					data <= x"7D48";
--				when '0' & x"5B" =>
--					data <= x"7D10";
--				when '0' & x"5C" =>
--					data <= x"7D0E";
--				when '0' & x"5D" =>
--					data <= x"9000";
--				when '0' & x"5E" =>
--					data <= x"910E";
--				when '0' & x"5F" =>
--					data <= x"911A";
--				when '0' & x"60" =>
--					data <= x"9131";
--				when '0' & x"61" =>
--					data <= x"915A";
--				when '0' & x"62" =>
--					data <= x"9169";
--				when '0' & x"63" =>
--					data <= x"9175";
--				when '0' & x"64" =>
--					data <= x"917E";
--				when '0' & x"65" =>
--					data <= x"9188";
--				when '0' & x"66" =>
--					data <= x"918F";
--				when '0' & x"67" =>
--					data <= x"9196";
--				when '0' & x"68" =>
--					data <= x"91A3";
--				when '0' & x"69" =>
--					data <= x"91AF";
--				when '0' & x"6A" =>
--					data <= x"91C4";
--				when '0' & x"6B" =>
--					data <= x"91D7";
--				when '0' & x"6C" =>
--					data <= x"91E8";
--				when '0' & x"6D" =>
--					data <= x"9120";
--				when '0' & x"6E" =>
--					data <= x"9200";
--				when '0' & x"6F" =>
--					data <= x"9306";
--				when '0' & x"70" =>
--					data <= x"93E3";
--				when '0' & x"71" =>
--					data <= x"9305";
--				when '0' & x"72" =>
--					data <= x"9305";
--				when '0' & x"73" =>
--					data <= x"9300";
--				when '0' & x"74" =>
--					data <= x"9600";
--				when '0' & x"75" =>
--					data <= x"9708";
--				when '0' & x"76" =>
--					data <= x"9719";
--				when '0' & x"77" =>
--					data <= x"9708";
--				when '0' & x"78" =>
--					data <= x"9719";
--				when '0' & x"79" =>
--					data <= x"9700";
--				when '0' & x"7A" =>
--					data <= x"C3ED";
--				when '0' & x"7B" =>
--					data <= x"A400";
--				when '0' & x"7C" =>
--					data <= x"A800";
--				when '0' & x"7D" =>
--					data <= x"C511";
--				when '0' & x"7E" =>
--					data <= x"C651";
--				when '0' & x"7F" =>
--					data <= x"BF80";
--				when '0' & x"80" =>
--					data <= x"C710";
--				when '0' & x"81" =>
--					data <= x"B666";
--				when '0' & x"82" =>
--					data <= x"B8A5";
--				when '0' & x"83" =>
--					data <= x"B764";
--				when '0' & x"84" =>
--					data <= x"B97C";
--				when '0' & x"85" =>
--					data <= x"B3AF";
--				when '0' & x"86" =>
--					data <= x"B497";
--				when '0' & x"87" =>
--					data <= x"B5FF";
--				when '0' & x"88" =>
--					data <= x"B0C5";
--				when '0' & x"89" =>
--					data <= x"B194";
--				when '0' & x"8A" =>
--					data <= x"B20F";
--				when '0' & x"8B" =>
--					data <= x"C45C";
--				when '0' & x"8C" =>
--					data <= x"C050";
--				when '0' & x"8D" =>
--					data <= x"C13C";
--				when '0' & x"8E" =>
--					data <= x"8C00";
--				when '0' & x"8F" =>
--					data <= x"863D";
--				when '0' & x"90" =>
--					data <= x"5000";
--				when '0' & x"91" =>
--					data <= x"51A0";
--				when '0' & x"92" =>
--					data <= x"5278";
--				when '0' & x"93" =>
--					data <= x"5300";
--				when '0' & x"94" =>
--					data <= x"5400";
--				when '0' & x"95" =>
--					data <= x"5500";
--				when '0' & x"96" =>
--					data <= x"5AA0";
--				when '0' & x"97" =>
--					data <= x"5B78";
--				when '0' & x"98" =>
--					data <= x"5C00";
--				when '0' & x"99" =>
--					data <= x"D382";
--				when '0' & x"9A" =>
--					data <= x"C3ED";
--				when '0' & x"9B" =>
--					data <= x"7F00";
--				when '0' & x"9C" =>
--					data <= x"DA08";
--				when '0' & x"9D" =>
--					data <= x"E51F";
--				when '0' & x"9E" =>
--					data <= x"E167";
--				when '0' & x"9F" =>
--					data <= x"E000";
--				when '0' & x"A0" =>
--					data <= x"DD7F";
--				when '0' & x"A1" =>
--					data <= x"0500";
--				when '0' & x"A2" =>
--					data <= x"FF01";
--				when '0' & x"A3" =>
--					data <= x"FF01";
--				when '0' & x"A4" =>
--					data <= x"FF01";
--				when '0' & x"A5" =>
--					data <= x"FF01";
--				when '0' & x"A6" =>
--					data <= x"FF01";
--				when '0' & x"A7" =>
--					data <= x"FF01";
--				when '0' & x"A8" =>
--					data <= x"FF01";
--				when '0' & x"A9" =>
--					data <= x"FF01";
--				when '0' & x"AA" =>
--					data <= x"FF01";
				when others =>
					data <= x"0000";
					finished <= '1';
					
				
				
				
				
				
				
				
				
				
--				when '0' & x"00" =>
--					data <= x"FF01";
--				when '0' & x"01" =>
--					data <= x"1100";
--				when '0' & x"02" =>
--					data <= x"1240";
--				when '0' & x"03" =>
--					data <= x"2A00";
--				when '0' & x"04" =>
--					data <= x"2B00";
--				when '0' & x"05" =>
--					data <= x"4600";
--				when '0' & x"06" =>
--					data <= x"4700";
--				when '0' & x"07" =>
--					data <= x"3D38";
--				when others =>
--					data <= x"0000";
--					finished <= '1';
					
					
					
					
					
				end case;
		end if;
	end process;

end INIT_RAM_ARCH;